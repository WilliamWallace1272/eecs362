module datapath (input clk, output [0:31] instruction);

    i_fetch I_FETCH(.clk(clk), .target()
    i_decode I_DECODE(.clk(clk), .



endmodule
